	
	
module simulator



//get result of what happened in one month
pub fn (mut sim Simulator) month_result_get(month int) ?{



}
