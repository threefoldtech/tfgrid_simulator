module tfgridsimulator

pub struct Node{
pub mut:
	nr_cu f32
	nr_su f32
}


